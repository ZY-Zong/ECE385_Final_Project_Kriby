module area1data (
	input  logic [17:0] addr,
	output logic [2:0] area1index
);
parameter[1:213839][2:0] data = {
	3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h0,3'h0,3'h7,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h7,3'h0,3'h0,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h6,3'h0,3'h5,3'h6,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h6,3'h0,3'h0,3'h5,3'h5,3'h6,3'h7,3'h0,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h5,3'h5,3'h6,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h5,3'h5,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h0,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h0,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h6,3'h6,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h2,3'h6,3'h6,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h6,3'h2,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h2,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h0,3'h0,3'h7,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h7,3'h0,3'h0,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h6,3'h0,3'h5,3'h6,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h6,3'h0,3'h0,3'h5,3'h5,3'h6,3'h7,3'h0,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h5,3'h5,3'h6,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h5,3'h5,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h1,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h1,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h0,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h6,3'h1,3'h5,3'h5,3'h1,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h5,3'h5,3'h1,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h6,3'h6,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h2,3'h1,3'h1,3'h5,3'h5,3'h5,3'h1,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h1,3'h1,3'h5,3'h5,3'h5,3'h1,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h1,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h1,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h1,3'h5,3'h5,3'h5,3'h5,3'h5,3'h1,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h1,3'h5,3'h5,3'h5,3'h5,3'h5,3'h1,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h1,3'h5,3'h5,3'h1,3'h1,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h5,3'h5,3'h1,3'h1,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h1,3'h5,3'h1,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h6,3'h5,3'h1,3'h5,3'h1,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h1,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h5,3'h5,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h5,3'h5,3'h2,3'h6,3'h5,3'h6,3'h1,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h0,3'h6,3'h1,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h5,3'h6,3'h6,3'h5,3'h5,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h0,3'h5,3'h5,3'h6,3'h6,3'h5,3'h6,3'h0,3'h6,3'h1,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h6,3'h0,3'h6,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h6,3'h5,3'h5,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h6,3'h6,3'h0,3'h6,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h0,3'h6,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h6,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h6,3'h6,3'h6,3'h0,3'h6,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h6,3'h5,3'h6,3'h2,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h7,3'h5,3'h7,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h5,3'h7,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h0,3'h4,3'h4,3'h4,3'h4,3'h4,3'h0,3'h0,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h0,3'h4,3'h4,3'h4,3'h4,3'h4,3'h0,3'h0,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h6,3'h7,3'h7,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h7,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h0,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h4,3'h4,3'h0,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h6,3'h6,3'h7,3'h7,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h7,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h0,3'h4,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h4,3'h7,3'h4,3'h4,3'h0,3'h4,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h4,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h7,3'h5,3'h7,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h5,3'h7,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h4,3'h4,3'h4,3'h4,3'h0,3'h0,3'h0,3'h0,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h4,3'h4,3'h4,3'h4,3'h0,3'h0,3'h0,3'h0,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h7,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h4,3'h4,3'h0,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h4,3'h4,3'h0,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h1,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h6,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h1,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h5,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h5,3'h5,3'h1,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h5,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h1,3'h1,3'h5,3'h5,3'h5,3'h1,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h6,3'h6,3'h6,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h1,3'h5,3'h5,3'h5,3'h5,3'h5,3'h1,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h1,3'h5,3'h5,3'h1,3'h1,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h1,3'h5,3'h1,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h7,3'h5,3'h5,3'h7,3'h5,3'h5,3'h6,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h7,3'h5,3'h5,3'h7,3'h5,3'h5,3'h6,3'h2,3'h2,3'h5,3'h5,3'h6,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h6,3'h1,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h5,3'h5,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h0,3'h5,3'h5,3'h5,3'h6,3'h5,3'h5,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h7,3'h7,3'h7,3'h5,3'h5,3'h6,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h7,3'h7,3'h7,3'h5,3'h5,3'h6,3'h2,3'h5,3'h5,3'h6,3'h5,3'h5,3'h5,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h0,3'h6,3'h1,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h5,3'h6,3'h6,3'h5,3'h5,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h0,3'h5,3'h5,3'h6,3'h6,3'h5,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h4,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h5,3'h6,3'h5,3'h6,3'h6,3'h5,3'h5,3'h0,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h0,3'h6,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h6,3'h5,3'h5,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h5,3'h5,3'h6,3'h6,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h7,3'h7,3'h7,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h4,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h7,3'h7,3'h7,3'h5,3'h5,3'h6,3'h6,3'h6,3'h5,3'h5,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h0,3'h6,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h6,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h0,3'h6,3'h6,3'h6,3'h5,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h7,3'h5,3'h5,3'h7,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h4,3'h6,3'h5,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h7,3'h5,3'h5,3'h7,3'h5,3'h5,3'h6,3'h6,3'h6,3'h0,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h6,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h7,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h4,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h7,3'h5,3'h5,3'h6,3'h6,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h1,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h5,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h4,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h4,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h5,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h4,3'h6,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h5,3'h7,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h6,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h7,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h6,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h7,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h6,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h5,3'h7,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h7,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h4,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h6,3'h4,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h4,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h6,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h6,3'h5,3'h0,3'h0,3'h5,3'h0,3'h5,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h6,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h6,3'h6,3'h6,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h6,3'h6,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h4,3'h6,3'h6,3'h6,3'h5,3'h0,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h4,3'h4,3'h4,3'h4,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h4,3'h4,3'h4,3'h4,3'h5,3'h5,3'h6,3'h6,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h6,3'h5,3'h5,3'h5,3'h0,3'h5,3'h0,3'h0,3'h5,3'h4,3'h4,3'h4,3'h4,3'h5,3'h5,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h6,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h6,3'h5,3'h5,3'h0,3'h0,3'h5,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h6,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h5,3'h0,3'h0,3'h5,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h5,3'h0,3'h0,3'h5,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h6,3'h6,3'h5,3'h5,3'h0,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h5,3'h0,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h5,3'h0,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h6,3'h6,3'h5,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h4,3'h6,3'h4,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h4,3'h4,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h4,3'h4,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h2,3'h2,3'h2,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h7,3'h7,3'h7,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h7,3'h7,3'h7,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h2,3'h2,3'h4,3'h4,3'h4,3'h4,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h7,3'h7,3'h7,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h4,3'h4,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h4,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h7,3'h7,3'h4,3'h7,3'h4,3'h4,3'h4,3'h4,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h4,3'h4,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h2,3'h4,3'h4,3'h7,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h2,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h4,3'h0,3'h0,3'h7,3'h7,3'h4,3'h7,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h4,3'h4,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h4,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h7,3'h4,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h4,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h4,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h4,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h4,3'h4,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h7,3'h7,3'h7,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h5,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h7,3'h7,3'h7,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h7,3'h7,3'h7,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h3,3'h7,3'h7,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h3,3'h3,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h7,3'h7,3'h7,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h7,3'h7,3'h7,3'h5,3'h1,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h5,3'h5,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h5,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h0,3'h0,3'h5,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h5,3'h1,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h7,3'h0,3'h5,3'h5,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h1,3'h1,3'h1,3'h5,3'h1,3'h1,3'h1,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h1,3'h5,3'h7,3'h7,3'h7,3'h1,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h7,3'h7,3'h3,3'h3,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h1,3'h5,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h5,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h3,3'h3,3'h3,3'h3,3'h3,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h5,3'h0,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h7,3'h7,3'h7,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0,3'h0
};
assign area1index = data[addr];
endmodule